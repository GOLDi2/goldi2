-------------------------------------------------------------------------------
-- Company:			Technische Universitaet Ilmenau
-- Engineer:		JP_CC <josepablo.chew@gmail.com>
--
-- Create Date:		30/04/2023
-- Design Name:		Warehouse sensor array
-- Module Name:		WH_SENSOR_ARRAY
-- Project Name:	GOLDi_FPGA_SRC
-- Target Devices:	LCMXO2-7000HC-4TG144C
-- Tool versions:	Lattice Diamond 3.12, Modelsim Lattice Edition,  
--
-- Dependencies:	-> GOLDI_COMM_STANDARD.vhd
--                  -> GOLDI_IO_STANDARD.vhd
--                  -> GOLDI_DATA_TYPES.vhd
--                  -> REGISTER_TABLE.vhd
--                  -> VIRTUAL_SENSOR_ARRAY.vhd
--
-- Revisions:
-- Revision V1.00.00 - File Created
-- Additional Comments: First commitment
-- 
-- Revision V2.00.00 - First release
-- Additional Comments:
--
-- Revision V4.00.00 - Module refactoring
-- Additional Comments: Change to the generic and port signal names to follow
--                      V4.00.00 naming convention. Correction of the 
--                      instantiated entities. Change to reset for the 
--                      virtual sensor arrays.
-------------------------------------------------------------------------------
--! Standard library
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--! Custom packages
library work;
use work.GOLDI_COMM_STANDARD.all;
use work.GOLDI_IO_STANDARD.all;
use work.GOLDI_DATA_TYPES.all;




--! @brief Possition sensor array for the GOLDi "Warehouse" Model
--! @details
--! The module consists of two sets of position values. 
--!
--! The first consists of the values gatherd from the physical switches accross the
--! model. These values are the limit sensors that prevent damage to the Warehouse.
--! Additionaly an inductive sensor indicates if the Warehouse crane is loaded. This
--! data is stored in the lowest register in the current 8-bit data system. (Data 
--! would be automatically strored in the lowest 8 bits if the data width is increased).
--!
--! The second group of values are "virtual" position values i.e. values calculated by
--! tracking the movement of the Warehouse crane using the x-axis and z-axis incremetal
--! encoders. The virtual sensors assert if the crane is located inside a given range
--! of the x or z axes. These values allow the use to allign the crane with one of the 
--! 50 loading bays before moving the content. The data generated by the virtual sensors
--! is stored in the upper 2 registers of the module. The 10 lowest bits [9:0] correspond
--! to the 10 x-axis sensors and the upper 5 [14:10] to the 5 z-axis sensors.
--!
--! | g_address	| Bit 7	| Bit 6 | Bit 5 | Bit 4 | Bit 3 | Bit 2 | Bit 1 | Bit 0 |
--! |----------:|:-----:|:- ---:|:-----:|:-----:|:-----:|:-----:|:-----:|:-----:|
--!	| +0		|       | ind   | z_pos | z_neg | y_pos | y_neg | z_pos | z_neg |
--! | +1        |           virtual_x_sensors [7:0]                      ||||||||
--! | +2        |       |virtual_z_sensors [14:10] |||||virutal_x_sensors [9:8]||
--! 
--! ***Lantency: 3cyc***
entity WH_SENSOR_ARRAY is
    generic(
        g_address           :   natural := 1;                                           --! Module's base address
        g_enc_x_invert      :   boolean := false;                                       --! Select x encoder positive direction [false -> CCW | true -> CC]
        g_enc_z_invert      :   boolean := false;                                       --! Select z encoder positive direction [false -> CCW | true -> CC]
        g_x_limit_sensors   :   sensor_limit_array(9 downto 0) := (others => (10,0));   --! X-axis loading bays position values (GOLDI_MODULE_CONFIG)
        g_z_limit_sensors   :   sensor_limit_array(4 downto 0) := (others => (10,0))    --! Z-axis loading bays position values (GOLDI_MODULE_CONFIG)
    );
    port(
        --General
        clk                 : in    std_logic;                                          --! System clock
        rst                 : in    std_logic;                                          --! Asynchronous reset
        ref_virtual_x       : in    std_logic;                                          --! Reset for x virtual sensor array
        ref_virtual_z       : in    std_logic;                                          --! Reset for z virtual sensor array
        --BUS slave interface
        sys_bus_i           : in    sbus_in;                                            --! BUS input signals [stb,we,adr,dat,tag]
        sys_bus_o           : out   sbus_out;                                           --! BUS output signals [dat,tag,mux]
        --Mechanical limit swiches
        p_lim_x_neg         : in    io_i;                                               --! X-Axis negative limit sensor
        p_lim_x_pos         : in    io_i;                                               --! X-Axis positive limit sensor
        p_lim_y_neg         : in    io_i;                                               --! Y-Axis negative limit sensor
        p_lim_y_pos         : in    io_i;                                               --! Y-Axis positive limit sensor
        p_lim_z_neg         : in    io_i;                                               --! Z-Axis negative limit sensor
        p_lim_z_pos         : in    io_i;                                               --! Z-Axis positive limit sensor
        p_inductive         : in    io_i;                                               --! Inductive sensor (active low)
        --Encoder signals
        p_channel_x_a       : in    io_i;                                               --! X-axis incremental encoder channel a
        p_channel_x_b       : in    io_i;                                               --! X-axis incremental encoder channel b
        p_channel_z_a       : in    io_i;                                               --! Z-axis incremental encoder channel a
        p_channel_z_b       : in    io_i                                                --! Z-axis incremental encoder channel b
    );
end entity WH_SENSOR_ARRAY;




--! General architecture
architecture RTL of WH_SENSOR_ARRAY is

    --****INTERNAL SIGNALS****
    --Memory
    constant memory_length  :   natural := getMemoryLength(23);
    constant reg_default    :   data_word_vector(memory_length-1 downto 0) := (others => (others => '0'));
    signal reg_data         :   data_word_vector(memory_length-1 downto 0); 
    --Virtual sensor reset
    signal rst_virtual_x    :   std_logic;
    signal rst_virtual_z    :   std_logic;
    --Sensor buffer
    signal sensor_buff      :   std_logic_vector(22 downto 0);


begin

    --****LIMIT SENSORS****
    -----------------------------------------------------------------------------------------------
    sensor_buff(0) <= p_lim_x_neg.dat;
    sensor_buff(1) <= p_lim_x_pos.dat;
    sensor_buff(2) <= p_lim_y_neg.dat;
    sensor_buff(3) <= p_lim_y_pos.dat;
    sensor_buff(4) <= p_lim_z_neg.dat;
    sensor_buff(5) <= p_lim_z_pos.dat;
    sensor_buff(6) <= not p_inductive.dat;
    sensor_buff(7) <= '0';
    -----------------------------------------------------------------------------------------------



    --****VIRTUAL SENSORS X AXIS****
    -----------------------------------------------------------------------------------------------
    rst_virtual_x <= rst or ref_virtual_x;

    X_SENSORS : entity work.VIRTUAL_SENSOR_ARRAY
    generic map(
        g_invert            => g_enc_x_invert,
        g_number_sensors    => 10,
        g_sensor_limits     => g_x_limit_sensors
    )
    port map(
        clk                 => clk,
        rst                 => rst_virtual_x,
        p_channel_a         => p_channel_x_a.dat,
        p_channel_b         => p_channel_x_b.dat,
        p_sensor_data       => sensor_buff(17 downto 8)
    );
    -----------------------------------------------------------------------------------------------



    --****VIRTUAL SENSORS Z AXIS****
    -----------------------------------------------------------------------------------------------
    rst_virtual_z <= rst or ref_virtual_z;
    
    Z_SENSORS : entity work.VIRTUAL_SENSOR_ARRAY
    generic map(
        g_invert            => g_enc_z_invert,
        g_number_sensors    => 5,
        g_sensor_limits     => g_z_limit_sensors
    )
    port map(
        clk                 => clk,
        rst                 => rst_virtual_z,
        p_channel_a         => p_channel_z_a.dat,
        p_channel_b         => p_channel_z_b.dat,
        p_sensor_data       => sensor_buff(22 downto 18)
    );
    -----------------------------------------------------------------------------------------------



    --****MEMORY****
    -----------------------------------------------------------------------------------------------
    MEMORY : entity work.REGISTER_TABLE
    generic map(
        g_address       => g_address,
        g_reg_number    => memory_length,
        g_def_values    => reg_default
    )
    port map(
        clk             => clk,
        rst             => rst,
        sys_bus_i       => sys_bus_i,
        sys_bus_o       => sys_bus_o,
        p_data_in       => reg_data,
        p_data_out      => open,
        p_read_stb      => open,
        p_write_stb     => open
    );
	
	reg_data <= setMemory(sensor_buff);
    -----------------------------------------------------------------------------------------------


end architecture; 
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package crossbar_config is
    constant config : work.crossbar.uconfig_word_vector(0 to 63) := (
        std_logic_vector(to_unsigned(0,8)),
        std_logic_vector(to_unsigned(1,8)),
        std_logic_vector(to_unsigned(2,8)),
        std_logic_vector(to_unsigned(3,8)),
        std_logic_vector(to_unsigned(4,8)),
        std_logic_vector(to_unsigned(5,8)),
        std_logic_vector(to_unsigned(6,8)),
        std_logic_vector(to_unsigned(7,8)),
        std_logic_vector(to_unsigned(8,8)),
        std_logic_vector(to_unsigned(9,8)),
        std_logic_vector(to_unsigned(10,8)),
        std_logic_vector(to_unsigned(11,8)),
        std_logic_vector(to_unsigned(12,8)),
        std_logic_vector(to_unsigned(13,8)),
        std_logic_vector(to_unsigned(14,8)),
        std_logic_vector(to_unsigned(15,8)),
        std_logic_vector(to_unsigned(16,8)),
        std_logic_vector(to_unsigned(17,8)),
        std_logic_vector(to_unsigned(18,8)),
        std_logic_vector(to_unsigned(19,8)),
        std_logic_vector(to_unsigned(20,8)),
        std_logic_vector(to_unsigned(21,8)),
        std_logic_vector(to_unsigned(22,8)),
        std_logic_vector(to_unsigned(23,8)),
        std_logic_vector(to_unsigned(24,8)),
        std_logic_vector(to_unsigned(25,8)),
        std_logic_vector(to_unsigned(26,8)),
        std_logic_vector(to_unsigned(27,8)),
        std_logic_vector(to_unsigned(28,8)),
        std_logic_vector(to_unsigned(29,8)),
        std_logic_vector(to_unsigned(30,8)),
        std_logic_vector(to_unsigned(31,8)),
        std_logic_vector(to_unsigned(32,8)),
        std_logic_vector(to_unsigned(33,8)),
        std_logic_vector(to_unsigned(34,8)),
        std_logic_vector(to_unsigned(35,8)),
        std_logic_vector(to_unsigned(36,8)),
        std_logic_vector(to_unsigned(37,8)),
        std_logic_vector(to_unsigned(38,8)),
        std_logic_vector(to_unsigned(39,8)),
        std_logic_vector(to_unsigned(40,8)),
        std_logic_vector(to_unsigned(41,8)),
        std_logic_vector(to_unsigned(42,8)),
        std_logic_vector(to_unsigned(43,8)),
        std_logic_vector(to_unsigned(44,8)),
        std_logic_vector(to_unsigned(45,8)),
        std_logic_vector(to_unsigned(46,8)),
        std_logic_vector(to_unsigned(47,8)),
        std_logic_vector(to_unsigned(48,8)),
        std_logic_vector(to_unsigned(49,8)),
        std_logic_vector(to_unsigned(50,8)),
        std_logic_vector(to_unsigned(51,8)),
        std_logic_vector(to_unsigned(52,8)),
        std_logic_vector(to_unsigned(53,8)),
        std_logic_vector(to_unsigned(54,8)),
        std_logic_vector(to_unsigned(55,8)),
        std_logic_vector(to_unsigned(56,8)),
        std_logic_vector(to_unsigned(57,8)),
        std_logic_vector(to_unsigned(58,8)),
        std_logic_vector(to_unsigned(59,8)),
        std_logic_vector(to_unsigned(60,8)),
        std_logic_vector(to_unsigned(61,8)),
        std_logic_vector(to_unsigned(62,8)),
        std_logic_vector(to_unsigned(63,8))
    );
end package crossbar_config;
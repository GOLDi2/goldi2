-------------------------------------------------------------------------------
-- Company:			Technische Universität Ilmenau
-- Engineer:		JP_CC <josepablo.chew@gmail.com>
--
-- Create Date:		15/04/2023
-- Design Name:		TMC2660 SPI Driver 
-- Module Name:		TMC2660_SPI
-- Project Name:	GOLDi_FPGA_SRC
-- Target Devices:	LCMXO2-7000HC-4TG144C
-- Tool versions:	Lattice Diamond 3.12, Modelsim Lattice Edition
--
-- Dependencies:    none
--
-- Revisions:
-- Revision V1.00.00 - File Created
-- Additional Comments: First commitment
--
-- Revision V2.00.00 - Default module version for release 1.00.00
-- Additional Comments: -  
-------------------------------------------------------------------------------
--! Use standard library
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;




--! @brief
--! @details
entity TMC2660_SPI is
    generic(
        CLOCK_FACTOR    :   natural := 8
    );
    port(
        --General
        clk             : in    std_logic;
        rst             : in    std_logic;
        --Parallel interface
        s_word_i_tready : out   std_logic;
        s_word_i_tvalid : in    std_logic;
        s_word_i_tdata  : in    std_logic_vector(19 downto 0);
        m_word_o_tvalid : out   std_logic;
        m_word_o_tdata  : out   std_logic_vector(19 downto 0);
        --Serial interface
        m_spi_sclk      : out   std_logic;
        m_spi_ncs       : out   std_logic;
        m_spi_mosi      : out   std_logic;
        m_spi_miso      : in    std_logic
    );
end entity TMC2660_SPI;




--! General architecture
architecture RTL of TMC2660_SPI is

    --****INTENAL SIGNALS****
    --Data buffers
    signal word_i_buff  :   std_logic_vector(19 downto 0);
    signal word_o_buff  :   std_logic_vector(19 downto 0);
    --Counters
    signal sclk_counter :   natural range 0 to CLOCK_FACTOR;
    signal bit_counter  :   natural range 0 to 19;
    --Flags
    signal s_ready_i    :   std_logic;
    signal m_valid_i    :   std_logic;
    signal tx_valid     :   std_logic;
    --State machine
    type spi_state is (IDLE, ENABLE, TRANSFER, DISABLE);
    signal spi_ps : spi_state := IDLE;


begin

    --****MODULE CONTROL****
    -----------------------------------------------------------------------------------------------
    STATE_MACHINE : process(clk)
    begin
        if(rising_edge(clk)) then
            
            --Control module parallel interface and spi transfer
            case spi_ps is
                when IDLE =>
                    word_i_buff <= s_word_i_tdata;
                    m_word_o_tdata <= word_o_buff;
                    --Start transfer once a new data word has been latched
                    if(s_word_i_tvalid = '1' and s_ready_i = '1') then
                        spi_ps <= ENABLE;
                    end if;

                when ENABLE =>
                    spi_ps <= TRANSFER;

                when TRANSFER =>
                    if(bit_counter = 19 and sclk_counter = CLOCK_FACTOR/2+1) then
                        spi_ps <= DISABLE;
                        tx_valid <= '1';
                    end if;

                when DISABLE =>
                    spi_ps <= IDLE;
                
            end case;

            
            --Reset module
            if(rst = '1') then
                word_i_buff <= (others => '0');
                tx_valid    <= '0';
                spi_ps      <= IDLE;
            end if;
        
        end if;
    end process;


    S_READY_FLAG_MANAGEMENT : process(spi_ps, tx_valid)
    begin
        --Manage ready flag
        if(spi_ps = IDLE) then
            s_ready_i <= '1';
        else
            s_ready_i <= '0';
        end if;
    end process;


    M_VALID_FLAG_MANAGEMENT : process(clk)
    begin
        if(rising_edge(clk)) then
            --Manage valid flag
            if(rst = '1') then
                m_valid_i <= '0';
            elsif(spi_ps = IDLE and tx_valid = '1') then
                m_valid_i <= '1';
            else
                m_valid_i <= '0';
            end if;
        end if;
    end process;

    s_word_i_tready <= s_ready_i;
    m_word_o_tvalid <= m_valid_i;
    -----------------------------------------------------------------------------------------------




    --****SPI INTERFACE****
    -----------------------------------------------------------------------------------------------
    SPI_SCLK_DIRVER : process(clk)
    begin
        if(rising_edge(clk)) then
            if(rst = '1') then
                m_spi_sclk <= '1';
            elsif(spi_ps /= TRANSFER) then
                m_spi_sclk <= '1';
            else
                if(sclk_counter < CLOCK_FACTOR/2) then
                    m_spi_sclk <= '0';
                else
                    m_spi_sclk <= '1';
                end if;
            end if;
        end if;
    end process;


    SPI_NCS_DRIVER : process(clk)
    begin
        if(rising_edge(clk)) then
            if(rst = '1') then
                m_spi_ncs <= '1';
            elsif(spi_ps = IDLE or spi_ps = DISABLE) then
                m_spi_ncs <= '1';
            else
                m_spi_ncs <= '0';
            end if;
        end if;
    end process;


    SPI_MOSI_DRIVER : process(clk)
    begin
        if(rising_edge(clk)) then
            if(rst = '1') then
                m_spi_mosi <= '0';
            elsif(spi_ps /= TRANSFER) then
                m_spi_mosi <= '0';
            else
                m_spi_mosi <= word_i_buff(19 - bit_counter);
            end if;
        end if;
    end process;


    SPI_MISO_DRIVER : process(clk)
    begin
        if(rising_edge(clk)) then
            if(rst = '1') then
                word_o_buff <= (others => '0');
            --Delay sample by two clk cycles to compensate for synchronizer delay
            elsif(spi_ps = TRANSFER and sclk_counter = CLOCK_FACTOR/2+1) then
                word_o_buff(19 - bit_counter) <= m_spi_miso; 
            end if;
        end if;
    end process;
    -----------------------------------------------------------------------------------------------




    --****COUNTERS****
    -----------------------------------------------------------------------------------------------
    SYSTEM_COUNTERS : process(clk)
    begin
        if(rising_edge(clk)) then
            if(rst = '1') then
                sclk_counter <= 0;
                bit_counter  <= 0;
            elsif(spi_ps /= TRANSFER) then
                sclk_counter <= 0;
                bit_counter  <= 0;
            else
                --Cycle a counter for serial clock signal
                if(sclk_counter = CLOCK_FACTOR-1) then
                    sclk_counter <= 0;
                else
                    sclk_counter <= sclk_counter + 1;
                end if;

                --Cycle a 20 counter for bit transfer
                if(bit_counter = 19 and sclk_counter = CLOCK_FACTOR-1) then
                    bit_counter <= 0;
                elsif(sclk_counter = CLOCK_FACTOR-1) then
                    bit_counter <= bit_counter + 1;
                end if;
            
            end if;
        end if;
    end process;
    -----------------------------------------------------------------------------------------------


end RTL;